package types is
    TYPE statetype IS (SB, S0, S1, S00, S01, S10, S11, RX, C, SUB, C2, SUM, TX);
end types;
